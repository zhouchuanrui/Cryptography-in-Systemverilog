//
//File: base_pkg.sv
//Device: 
//Created:  2017-4-9 15:32:20
//Description: base package
//Revisions: 
//2017-4-9 15:32:29: created
//

`ifndef __BASE_PKG
`define __BASE_PKG
package base_pkg;

    `include "base_macros.svh"
    `include "LogBase.svh"
endpackage
`endif

