//
//File: test_pkg.sv
//Device: 
//Created:  2017-4-18 22:55:14
//Description: test package
//Revisions: 
//2017-4-18 22:55:25: created
//

package test_pkg;
    `include "base_macros.svh"
    import base_pkg::LogBase;

    `include "TestFactory.svh"

    `include "demo_test.svh"

    `include "aes_test.svh"
    `include "des_test.svh"
    `include "tdea_test.svh"
endpackage

